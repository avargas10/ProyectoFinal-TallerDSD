`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   18:10:04 11/27/2017
// Design Name:   topLevelModule
// Module Name:   C:/Users/Andres Vargas/Documents/Verilog Projects/microProcessor/microProcessor/total_test.v
// Project Name:  microProcessor
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: topLevelModule
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module total_test;

	// Inputs
	reg clk;
	reg reset;

	// Outputs
	wire [31:0] WriteData,DataAdr;
	wire MemWrite;
	// Instantiate the Unit Under Test (UUT)
	topLevelModule uut (
		.clk(clk), 
		.reset(reset),
		.WriteData(WriteData),
		.DataAdr(DataAdr),
		.MemWrite(MemWrite)		
	);

	initial
		begin
			reset <= 1; # 22; reset <= 0;
		end
// generate clock to sequence tests
always
	begin
		clk <= 1; # 5; clk <= 0; # 5;
	end
	
// check that 7 gets written to address 0x64
// at end of program
always @(negedge clk)
		begin
		if(MemWrite) begin
			if(DataAdr === 100 & WriteData === 7) begin
					$display("Simulation succeeded");
					$stop;
				end else if (DataAdr !== 96) begin
					$display("Simulation failed");
					$stop;
				end
			end
		end
endmodule

